library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;
library work;
use work.Common.all;

entity Sigmoid is
port (
	arg 	: in fixed_point;
	ret 	: out fixed_point
);
end Sigmoid;

architecture Behavioral of Sigmoid is
	begin
	process (arg) is
	begin
		if arg < -4096 then
			ret <= to_fixed_point(0);
		elsif arg > 4096 then
			ret <= to_fixed_point(1024);
		elsif arg > to_fixed_point(-4096) and arg <= to_fixed_point(-4096) then
			ret <= to_fixed_point(18);
		elsif arg > to_fixed_point(-4096) and arg <= to_fixed_point(-4044) then
			ret <= to_fixed_point(19);
		elsif arg > to_fixed_point(-4044) and arg <= to_fixed_point(-3993) then
			ret <= to_fixed_point(20);
		elsif arg > to_fixed_point(-3993) and arg <= to_fixed_point(-3942) then
			ret <= to_fixed_point(21);
		elsif arg > to_fixed_point(-3942) and arg <= to_fixed_point(-3891) then
			ret <= to_fixed_point(22);
		elsif arg > to_fixed_point(-3891) and arg <= to_fixed_point(-3840) then
			ret <= to_fixed_point(24);
		elsif arg > to_fixed_point(-3840) and arg <= to_fixed_point(-3788) then
			ret <= to_fixed_point(25);
		elsif arg > to_fixed_point(-3788) and arg <= to_fixed_point(-3737) then
			ret <= to_fixed_point(26);
		elsif arg > to_fixed_point(-3737) and arg <= to_fixed_point(-3686) then
			ret <= to_fixed_point(27);
		elsif arg > to_fixed_point(-3686) and arg <= to_fixed_point(-3635) then
			ret <= to_fixed_point(29);
		elsif arg > to_fixed_point(-3635) and arg <= to_fixed_point(-3584) then
			ret <= to_fixed_point(30);
		elsif arg > to_fixed_point(-3584) and arg <= to_fixed_point(-3532) then
			ret <= to_fixed_point(32);
		elsif arg > to_fixed_point(-3532) and arg <= to_fixed_point(-3481) then
			ret <= to_fixed_point(33);
		elsif arg > to_fixed_point(-3481) and arg <= to_fixed_point(-3430) then
			ret <= to_fixed_point(35);
		elsif arg > to_fixed_point(-3430) and arg <= to_fixed_point(-3379) then
			ret <= to_fixed_point(36);
		elsif arg > to_fixed_point(-3379) and arg <= to_fixed_point(-3328) then
			ret <= to_fixed_point(38);
		elsif arg > to_fixed_point(-3328) and arg <= to_fixed_point(-3276) then
			ret <= to_fixed_point(40);
		elsif arg > to_fixed_point(-3276) and arg <= to_fixed_point(-3225) then
			ret <= to_fixed_point(42);
		elsif arg > to_fixed_point(-3225) and arg <= to_fixed_point(-3174) then
			ret <= to_fixed_point(44);
		elsif arg > to_fixed_point(-3174) and arg <= to_fixed_point(-3123) then
			ret <= to_fixed_point(46);
		elsif arg > to_fixed_point(-3123) and arg <= to_fixed_point(-3072) then
			ret <= to_fixed_point(49);
		elsif arg > to_fixed_point(-3072) and arg <= to_fixed_point(-3020) then
			ret <= to_fixed_point(51);
		elsif arg > to_fixed_point(-3020) and arg <= to_fixed_point(-2969) then
			ret <= to_fixed_point(53);
		elsif arg > to_fixed_point(-2969) and arg <= to_fixed_point(-2918) then
			ret <= to_fixed_point(56);
		elsif arg > to_fixed_point(-2918) and arg <= to_fixed_point(-2867) then
			ret <= to_fixed_point(59);
		elsif arg > to_fixed_point(-2867) and arg <= to_fixed_point(-2816) then
			ret <= to_fixed_point(62);
		elsif arg > to_fixed_point(-2816) and arg <= to_fixed_point(-2764) then
			ret <= to_fixed_point(65);
		elsif arg > to_fixed_point(-2764) and arg <= to_fixed_point(-2713) then
			ret <= to_fixed_point(68);
		elsif arg > to_fixed_point(-2713) and arg <= to_fixed_point(-2662) then
			ret <= to_fixed_point(71);
		elsif arg > to_fixed_point(-2662) and arg <= to_fixed_point(-2611) then
			ret <= to_fixed_point(74);
		elsif arg > to_fixed_point(-2611) and arg <= to_fixed_point(-2560) then
			ret <= to_fixed_point(78);
		elsif arg > to_fixed_point(-2560) and arg <= to_fixed_point(-2508) then
			ret <= to_fixed_point(81);
		elsif arg > to_fixed_point(-2508) and arg <= to_fixed_point(-2457) then
			ret <= to_fixed_point(85);
		elsif arg > to_fixed_point(-2457) and arg <= to_fixed_point(-2406) then
			ret <= to_fixed_point(89);
		elsif arg > to_fixed_point(-2406) and arg <= to_fixed_point(-2355) then
			ret <= to_fixed_point(93);
		elsif arg > to_fixed_point(-2355) and arg <= to_fixed_point(-2304) then
			ret <= to_fixed_point(98);
		elsif arg > to_fixed_point(-2304) and arg <= to_fixed_point(-2252) then
			ret <= to_fixed_point(102);
		elsif arg > to_fixed_point(-2252) and arg <= to_fixed_point(-2201) then
			ret <= to_fixed_point(107);
		elsif arg > to_fixed_point(-2201) and arg <= to_fixed_point(-2150) then
			ret <= to_fixed_point(112);
		elsif arg > to_fixed_point(-2150) and arg <= to_fixed_point(-2099) then
			ret <= to_fixed_point(117);
		elsif arg > to_fixed_point(-2099) and arg <= to_fixed_point(-2048) then
			ret <= to_fixed_point(122);
		elsif arg > to_fixed_point(-2048) and arg <= to_fixed_point(-1996) then
			ret <= to_fixed_point(128);
		elsif arg > to_fixed_point(-1996) and arg <= to_fixed_point(-1945) then
			ret <= to_fixed_point(133);
		elsif arg > to_fixed_point(-1945) and arg <= to_fixed_point(-1894) then
			ret <= to_fixed_point(139);
		elsif arg > to_fixed_point(-1894) and arg <= to_fixed_point(-1843) then
			ret <= to_fixed_point(145);
		elsif arg > to_fixed_point(-1843) and arg <= to_fixed_point(-1792) then
			ret <= to_fixed_point(152);
		elsif arg > to_fixed_point(-1792) and arg <= to_fixed_point(-1740) then
			ret <= to_fixed_point(158);
		elsif arg > to_fixed_point(-1740) and arg <= to_fixed_point(-1689) then
			ret <= to_fixed_point(165);
		elsif arg > to_fixed_point(-1689) and arg <= to_fixed_point(-1638) then
			ret <= to_fixed_point(172);
		elsif arg > to_fixed_point(-1638) and arg <= to_fixed_point(-1587) then
			ret <= to_fixed_point(179);
		elsif arg > to_fixed_point(-1587) and arg <= to_fixed_point(-1536) then
			ret <= to_fixed_point(187);
		elsif arg > to_fixed_point(-1536) and arg <= to_fixed_point(-1484) then
			ret <= to_fixed_point(195);
		elsif arg > to_fixed_point(-1484) and arg <= to_fixed_point(-1433) then
			ret <= to_fixed_point(203);
		elsif arg > to_fixed_point(-1433) and arg <= to_fixed_point(-1382) then
			ret <= to_fixed_point(211);
		elsif arg > to_fixed_point(-1382) and arg <= to_fixed_point(-1331) then
			ret <= to_fixed_point(219);
		elsif arg > to_fixed_point(-1331) and arg <= to_fixed_point(-1280) then
			ret <= to_fixed_point(228);
		elsif arg > to_fixed_point(-1280) and arg <= to_fixed_point(-1228) then
			ret <= to_fixed_point(237);
		elsif arg > to_fixed_point(-1228) and arg <= to_fixed_point(-1177) then
			ret <= to_fixed_point(246);
		elsif arg > to_fixed_point(-1177) and arg <= to_fixed_point(-1126) then
			ret <= to_fixed_point(256);
		elsif arg > to_fixed_point(-1126) and arg <= to_fixed_point(-1075) then
			ret <= to_fixed_point(265);
		elsif arg > to_fixed_point(-1075) and arg <= to_fixed_point(-1024) then
			ret <= to_fixed_point(275);
		elsif arg > to_fixed_point(-1024) and arg <= to_fixed_point(-972) then
			ret <= to_fixed_point(286);
		elsif arg > to_fixed_point(-972) and arg <= to_fixed_point(-921) then
			ret <= to_fixed_point(296);
		elsif arg > to_fixed_point(-921) and arg <= to_fixed_point(-870) then
			ret <= to_fixed_point(307);
		elsif arg > to_fixed_point(-870) and arg <= to_fixed_point(-819) then
			ret <= to_fixed_point(318);
		elsif arg > to_fixed_point(-819) and arg <= to_fixed_point(-768) then
			ret <= to_fixed_point(329);
		elsif arg > to_fixed_point(-768) and arg <= to_fixed_point(-716) then
			ret <= to_fixed_point(340);
		elsif arg > to_fixed_point(-716) and arg <= to_fixed_point(-665) then
			ret <= to_fixed_point(351);
		elsif arg > to_fixed_point(-665) and arg <= to_fixed_point(-614) then
			ret <= to_fixed_point(363);
		elsif arg > to_fixed_point(-614) and arg <= to_fixed_point(-563) then
			ret <= to_fixed_point(375);
		elsif arg > to_fixed_point(-563) and arg <= to_fixed_point(-512) then
			ret <= to_fixed_point(387);
		elsif arg > to_fixed_point(-512) and arg <= to_fixed_point(-460) then
			ret <= to_fixed_point(399);
		elsif arg > to_fixed_point(-460) and arg <= to_fixed_point(-409) then
			ret <= to_fixed_point(411);
		elsif arg > to_fixed_point(-409) and arg <= to_fixed_point(-358) then
			ret <= to_fixed_point(423);
		elsif arg > to_fixed_point(-358) and arg <= to_fixed_point(-307) then
			ret <= to_fixed_point(436);
		elsif arg > to_fixed_point(-307) and arg <= to_fixed_point(-256) then
			ret <= to_fixed_point(448);
		elsif arg > to_fixed_point(-256) and arg <= to_fixed_point(-204) then
			ret <= to_fixed_point(461);
		elsif arg > to_fixed_point(-204) and arg <= to_fixed_point(-153) then
			ret <= to_fixed_point(474);
		elsif arg > to_fixed_point(-153) and arg <= to_fixed_point(-102) then
			ret <= to_fixed_point(487);
		elsif arg > to_fixed_point(-102) and arg <= to_fixed_point(-51) then
			ret <= to_fixed_point(499);
		elsif arg > to_fixed_point(-51) and arg <= to_fixed_point(0) then
			ret <= to_fixed_point(512);
		elsif arg > to_fixed_point(0) and arg <= to_fixed_point(51) then
			ret <= to_fixed_point(525);
		elsif arg > to_fixed_point(51) and arg <= to_fixed_point(102) then
			ret <= to_fixed_point(537);
		elsif arg > to_fixed_point(102) and arg <= to_fixed_point(153) then
			ret <= to_fixed_point(550);
		elsif arg > to_fixed_point(153) and arg <= to_fixed_point(204) then
			ret <= to_fixed_point(563);
		elsif arg > to_fixed_point(204) and arg <= to_fixed_point(256) then
			ret <= to_fixed_point(576);
		elsif arg > to_fixed_point(256) and arg <= to_fixed_point(307) then
			ret <= to_fixed_point(588);
		elsif arg > to_fixed_point(307) and arg <= to_fixed_point(358) then
			ret <= to_fixed_point(601);
		elsif arg > to_fixed_point(358) and arg <= to_fixed_point(409) then
			ret <= to_fixed_point(613);
		elsif arg > to_fixed_point(409) and arg <= to_fixed_point(460) then
			ret <= to_fixed_point(625);
		elsif arg > to_fixed_point(460) and arg <= to_fixed_point(512) then
			ret <= to_fixed_point(637);
		elsif arg > to_fixed_point(512) and arg <= to_fixed_point(563) then
			ret <= to_fixed_point(649);
		elsif arg > to_fixed_point(563) and arg <= to_fixed_point(614) then
			ret <= to_fixed_point(661);
		elsif arg > to_fixed_point(614) and arg <= to_fixed_point(665) then
			ret <= to_fixed_point(673);
		elsif arg > to_fixed_point(665) and arg <= to_fixed_point(716) then
			ret <= to_fixed_point(684);
		elsif arg > to_fixed_point(716) and arg <= to_fixed_point(768) then
			ret <= to_fixed_point(695);
		elsif arg > to_fixed_point(768) and arg <= to_fixed_point(819) then
			ret <= to_fixed_point(706);
		elsif arg > to_fixed_point(819) and arg <= to_fixed_point(870) then
			ret <= to_fixed_point(717);
		elsif arg > to_fixed_point(870) and arg <= to_fixed_point(921) then
			ret <= to_fixed_point(728);
		elsif arg > to_fixed_point(921) and arg <= to_fixed_point(972) then
			ret <= to_fixed_point(738);
		elsif arg > to_fixed_point(972) and arg <= to_fixed_point(1024) then
			ret <= to_fixed_point(749);
		elsif arg > to_fixed_point(1024) and arg <= to_fixed_point(1075) then
			ret <= to_fixed_point(759);
		elsif arg > to_fixed_point(1075) and arg <= to_fixed_point(1126) then
			ret <= to_fixed_point(768);
		elsif arg > to_fixed_point(1126) and arg <= to_fixed_point(1177) then
			ret <= to_fixed_point(778);
		elsif arg > to_fixed_point(1177) and arg <= to_fixed_point(1228) then
			ret <= to_fixed_point(787);
		elsif arg > to_fixed_point(1228) and arg <= to_fixed_point(1280) then
			ret <= to_fixed_point(796);
		elsif arg > to_fixed_point(1280) and arg <= to_fixed_point(1331) then
			ret <= to_fixed_point(805);
		elsif arg > to_fixed_point(1331) and arg <= to_fixed_point(1382) then
			ret <= to_fixed_point(813);
		elsif arg > to_fixed_point(1382) and arg <= to_fixed_point(1433) then
			ret <= to_fixed_point(821);
		elsif arg > to_fixed_point(1433) and arg <= to_fixed_point(1484) then
			ret <= to_fixed_point(829);
		elsif arg > to_fixed_point(1484) and arg <= to_fixed_point(1536) then
			ret <= to_fixed_point(837);
		elsif arg > to_fixed_point(1536) and arg <= to_fixed_point(1587) then
			ret <= to_fixed_point(845);
		elsif arg > to_fixed_point(1587) and arg <= to_fixed_point(1638) then
			ret <= to_fixed_point(852);
		elsif arg > to_fixed_point(1638) and arg <= to_fixed_point(1689) then
			ret <= to_fixed_point(859);
		elsif arg > to_fixed_point(1689) and arg <= to_fixed_point(1740) then
			ret <= to_fixed_point(866);
		elsif arg > to_fixed_point(1740) and arg <= to_fixed_point(1792) then
			ret <= to_fixed_point(872);
		elsif arg > to_fixed_point(1792) and arg <= to_fixed_point(1843) then
			ret <= to_fixed_point(879);
		elsif arg > to_fixed_point(1843) and arg <= to_fixed_point(1894) then
			ret <= to_fixed_point(885);
		elsif arg > to_fixed_point(1894) and arg <= to_fixed_point(1945) then
			ret <= to_fixed_point(891);
		elsif arg > to_fixed_point(1945) and arg <= to_fixed_point(1996) then
			ret <= to_fixed_point(896);
		elsif arg > to_fixed_point(1996) and arg <= to_fixed_point(2048) then
			ret <= to_fixed_point(902);
		elsif arg > to_fixed_point(2048) and arg <= to_fixed_point(2099) then
			ret <= to_fixed_point(907);
		elsif arg > to_fixed_point(2099) and arg <= to_fixed_point(2150) then
			ret <= to_fixed_point(912);
		elsif arg > to_fixed_point(2150) and arg <= to_fixed_point(2201) then
			ret <= to_fixed_point(917);
		elsif arg > to_fixed_point(2201) and arg <= to_fixed_point(2252) then
			ret <= to_fixed_point(922);
		elsif arg > to_fixed_point(2252) and arg <= to_fixed_point(2304) then
			ret <= to_fixed_point(926);
		elsif arg > to_fixed_point(2304) and arg <= to_fixed_point(2355) then
			ret <= to_fixed_point(931);
		elsif arg > to_fixed_point(2355) and arg <= to_fixed_point(2406) then
			ret <= to_fixed_point(935);
		elsif arg > to_fixed_point(2406) and arg <= to_fixed_point(2457) then
			ret <= to_fixed_point(939);
		elsif arg > to_fixed_point(2457) and arg <= to_fixed_point(2508) then
			ret <= to_fixed_point(943);
		elsif arg > to_fixed_point(2508) and arg <= to_fixed_point(2560) then
			ret <= to_fixed_point(946);
		elsif arg > to_fixed_point(2560) and arg <= to_fixed_point(2611) then
			ret <= to_fixed_point(950);
		elsif arg > to_fixed_point(2611) and arg <= to_fixed_point(2662) then
			ret <= to_fixed_point(953);
		elsif arg > to_fixed_point(2662) and arg <= to_fixed_point(2713) then
			ret <= to_fixed_point(956);
		elsif arg > to_fixed_point(2713) and arg <= to_fixed_point(2764) then
			ret <= to_fixed_point(959);
		elsif arg > to_fixed_point(2764) and arg <= to_fixed_point(2816) then
			ret <= to_fixed_point(962);
		elsif arg > to_fixed_point(2816) and arg <= to_fixed_point(2867) then
			ret <= to_fixed_point(965);
		elsif arg > to_fixed_point(2867) and arg <= to_fixed_point(2918) then
			ret <= to_fixed_point(968);
		elsif arg > to_fixed_point(2918) and arg <= to_fixed_point(2969) then
			ret <= to_fixed_point(971);
		elsif arg > to_fixed_point(2969) and arg <= to_fixed_point(3020) then
			ret <= to_fixed_point(973);
		elsif arg > to_fixed_point(3020) and arg <= to_fixed_point(3072) then
			ret <= to_fixed_point(975);
		elsif arg > to_fixed_point(3072) and arg <= to_fixed_point(3123) then
			ret <= to_fixed_point(978);
		elsif arg > to_fixed_point(3123) and arg <= to_fixed_point(3174) then
			ret <= to_fixed_point(980);
		elsif arg > to_fixed_point(3174) and arg <= to_fixed_point(3225) then
			ret <= to_fixed_point(982);
		elsif arg > to_fixed_point(3225) and arg <= to_fixed_point(3276) then
			ret <= to_fixed_point(984);
		elsif arg > to_fixed_point(3276) and arg <= to_fixed_point(3328) then
			ret <= to_fixed_point(986);
		elsif arg > to_fixed_point(3328) and arg <= to_fixed_point(3379) then
			ret <= to_fixed_point(988);
		elsif arg > to_fixed_point(3379) and arg <= to_fixed_point(3430) then
			ret <= to_fixed_point(989);
		elsif arg > to_fixed_point(3430) and arg <= to_fixed_point(3481) then
			ret <= to_fixed_point(991);
		elsif arg > to_fixed_point(3481) and arg <= to_fixed_point(3532) then
			ret <= to_fixed_point(992);
		elsif arg > to_fixed_point(3532) and arg <= to_fixed_point(3584) then
			ret <= to_fixed_point(994);
		elsif arg > to_fixed_point(3584) and arg <= to_fixed_point(3635) then
			ret <= to_fixed_point(995);
		elsif arg > to_fixed_point(3635) and arg <= to_fixed_point(3686) then
			ret <= to_fixed_point(997);
		elsif arg > to_fixed_point(3686) and arg <= to_fixed_point(3737) then
			ret <= to_fixed_point(998);
		elsif arg > to_fixed_point(3737) and arg <= to_fixed_point(3788) then
			ret <= to_fixed_point(999);
		elsif arg > to_fixed_point(3788) and arg <= to_fixed_point(3840) then
			ret <= to_fixed_point(1000);
		elsif arg > to_fixed_point(3840) and arg <= to_fixed_point(3891) then
			ret <= to_fixed_point(1002);
		elsif arg > to_fixed_point(3891) and arg <= to_fixed_point(3942) then
			ret <= to_fixed_point(1003);
		elsif arg > to_fixed_point(3942) and arg <= to_fixed_point(3993) then
			ret <= to_fixed_point(1004);
		elsif arg > to_fixed_point(3993) and arg <= to_fixed_point(4044) then
			ret <= to_fixed_point(1005);
		elsif arg > to_fixed_point(4044) and arg <= to_fixed_point(4044) then
			ret <= to_fixed_point(1005);
		else
			ret <= factor;
		end if;
	end process;
end Behavioral;
